magic
tech scmos
timestamp 1731229290
<< nwell >>
rect -17 -32 191 38
<< polysilicon >>
rect 5 13 7 21
rect 44 13 46 17
rect 75 9 80 14
rect 111 13 113 18
rect 152 13 154 19
rect 5 -16 7 -11
rect 44 -16 46 -11
rect 75 -16 80 -11
rect 111 -20 113 -11
rect 152 -14 154 -11
rect 8 -45 10 -38
rect 47 -43 49 -36
rect 80 -43 82 -36
rect 120 -43 122 -36
rect 8 -57 10 -50
rect 47 -61 49 -53
rect 80 -60 82 -53
rect 120 -56 122 -53
rect 47 -81 49 -78
rect 80 -81 82 -74
rect 120 -81 122 -78
rect 47 -106 49 -91
rect 80 -98 82 -91
rect 120 -94 122 -91
<< ndiffusion >>
rect 5 -50 8 -45
rect 10 -50 13 -45
rect 44 -53 47 -43
rect 49 -53 52 -43
rect 77 -53 80 -43
rect 82 -53 85 -43
rect 117 -53 120 -43
rect 122 -53 125 -43
rect 44 -91 47 -81
rect 49 -91 52 -81
rect 77 -91 80 -81
rect 82 -91 85 -81
rect 117 -91 120 -81
rect 122 -91 125 -81
<< pdiffusion >>
rect 0 9 5 13
rect -4 -11 5 9
rect 7 -7 17 13
rect 7 -11 13 -7
rect 39 9 44 13
rect 35 -11 44 9
rect 46 -7 56 13
rect 106 9 111 13
rect 46 -11 52 -7
rect 71 5 75 9
rect 67 -11 75 5
rect 80 -7 89 9
rect 80 -11 85 -7
rect 102 -11 111 9
rect 113 -7 123 13
rect 113 -11 119 -7
rect 147 9 152 13
rect 143 -11 152 9
rect 154 -7 164 13
rect 154 -11 160 -7
<< metal1 >>
rect -8 31 -4 35
rect 0 31 5 35
rect 9 31 14 35
rect 18 31 23 35
rect 27 31 32 35
rect 36 31 41 35
rect 45 31 50 35
rect 54 31 58 35
rect 62 31 67 35
rect 71 31 76 35
rect 80 31 85 35
rect 89 31 94 35
rect 98 31 102 35
rect 106 31 110 35
rect 114 31 118 35
rect 122 31 126 35
rect 130 31 135 35
rect 139 31 143 35
rect 147 31 151 35
rect 155 31 161 35
rect 165 31 169 35
rect 173 31 175 35
rect -4 13 0 31
rect 11 17 27 21
rect -7 -16 1 -12
rect 13 -32 17 -11
rect 23 -12 27 17
rect 35 13 39 31
rect 67 9 71 31
rect 102 21 133 25
rect 102 13 106 21
rect 117 14 119 18
rect 23 -16 40 -12
rect 4 -36 17 -32
rect 52 -32 56 -11
rect 85 -16 89 -11
rect 79 -20 107 -16
rect 4 -38 8 -36
rect 13 -45 17 -36
rect 23 -40 43 -36
rect 1 -114 5 -50
rect 23 -53 27 -40
rect 52 -43 56 -36
rect 14 -57 27 -53
rect 65 -40 76 -36
rect 40 -68 44 -53
rect 65 -57 69 -40
rect 85 -43 89 -20
rect 119 -26 123 -11
rect 129 -16 133 21
rect 143 13 147 31
rect 158 15 180 19
rect 160 -16 164 -11
rect 129 -20 164 -16
rect 176 -26 180 15
rect 119 -30 180 -26
rect 53 -61 69 -57
rect 103 -40 116 -36
rect 73 -65 77 -53
rect 103 -56 107 -40
rect 125 -43 129 -30
rect 86 -60 107 -56
rect 40 -72 56 -68
rect 73 -69 89 -65
rect 52 -81 56 -72
rect 65 -78 76 -74
rect 40 -114 44 -91
rect 65 -102 69 -78
rect 85 -81 89 -69
rect 113 -66 117 -53
rect 113 -70 129 -66
rect 53 -106 69 -102
rect 104 -78 118 -74
rect 73 -114 77 -91
rect 104 -94 108 -78
rect 125 -81 129 -70
rect 86 -98 108 -94
rect 113 -114 117 -91
rect 4 -118 8 -114
rect 12 -118 16 -114
rect 20 -118 25 -114
rect 29 -118 34 -114
rect 38 -118 43 -114
rect 47 -118 53 -114
rect 57 -118 63 -114
rect 67 -118 72 -114
rect 76 -118 81 -114
rect 85 -118 89 -114
rect 93 -118 98 -114
rect 102 -118 107 -114
rect 111 -118 116 -114
rect 120 -118 125 -114
rect 129 -118 134 -114
rect 138 -118 142 -114
<< metal2 >>
rect 56 -36 62 -32
rect 58 -94 62 -36
rect 53 -98 62 -94
<< ntransistor >>
rect 8 -50 10 -45
rect 47 -53 49 -43
rect 80 -53 82 -43
rect 120 -53 122 -43
rect 47 -91 49 -81
rect 80 -91 82 -81
rect 120 -91 122 -81
<< ptransistor >>
rect 5 -11 7 13
rect 44 -11 46 13
rect 75 -11 80 9
rect 111 -11 113 13
rect 152 -11 154 13
<< polycontact >>
rect 7 17 11 21
rect 113 14 117 18
rect 154 15 158 19
rect 1 -16 5 -12
rect 40 -16 44 -12
rect 75 -20 79 -16
rect 107 -20 111 -16
rect 4 -42 8 -38
rect 43 -40 47 -36
rect 76 -40 80 -36
rect 116 -40 120 -36
rect 10 -57 14 -53
rect 49 -61 53 -57
rect 82 -60 86 -56
rect 76 -78 80 -74
rect 118 -78 122 -74
rect 49 -98 53 -94
rect 82 -98 86 -94
rect 49 -106 53 -102
<< ndcontact >>
rect 1 -50 5 -45
rect 13 -50 17 -45
rect 40 -53 44 -43
rect 52 -53 56 -43
rect 73 -53 77 -43
rect 85 -53 89 -43
rect 113 -53 117 -43
rect 125 -53 129 -43
rect 40 -91 44 -81
rect 52 -91 56 -81
rect 73 -91 77 -81
rect 85 -91 89 -81
rect 113 -91 117 -81
rect 125 -91 129 -81
<< pdcontact >>
rect -4 9 0 13
rect 13 -11 17 -7
rect 35 9 39 13
rect 102 9 106 13
rect 52 -11 56 -7
rect 67 5 71 9
rect 85 -11 89 -7
rect 119 -11 123 -7
rect 143 9 147 13
rect 160 -11 164 -7
<< m2contact >>
rect 52 -36 56 -32
<< psubstratepcontact >>
rect 0 -118 4 -114
rect 8 -118 12 -114
rect 16 -118 20 -114
rect 25 -118 29 -114
rect 34 -118 38 -114
rect 43 -118 47 -114
rect 53 -118 57 -114
rect 63 -118 67 -114
rect 72 -118 76 -114
rect 81 -118 85 -114
rect 89 -118 93 -114
rect 98 -118 102 -114
rect 107 -118 111 -114
rect 116 -118 120 -114
rect 125 -118 129 -114
rect 134 -118 138 -114
<< nsubstratencontact >>
rect -12 31 -8 35
rect -4 31 0 35
rect 5 31 9 35
rect 14 31 18 35
rect 23 31 27 35
rect 32 31 36 35
rect 41 31 45 35
rect 50 31 54 35
rect 58 31 62 35
rect 67 31 71 35
rect 76 31 80 35
rect 85 31 89 35
rect 94 31 98 35
rect 102 31 106 35
rect 110 31 114 35
rect 118 31 122 35
rect 126 31 130 35
rect 135 31 139 35
rect 143 31 147 35
rect 151 31 155 35
rect 161 31 165 35
rect 169 31 173 35
<< labels >>
rlabel metal1 70 -116 70 -116 1 gnd
rlabel metal1 -7 -16 -7 -12 1 vbiasp
rlabel metal1 119 14 119 18 1 vbias2
rlabel metal1 54 -106 54 -102 1 vbias4
rlabel metal1 160 15 160 19 1 vbias1
rlabel metal1 55 -61 55 -57 1 vbias3
rlabel metal1 81 33 81 33 5 vdd
<< end >>
