magic
tech scmos
timestamp 1731145861
<< nwell >>
rect -33 -59 32 51
<< polysilicon >>
rect -1 30 1 33
rect -1 5 1 6
rect -1 -27 1 -24
rect -1 -52 1 -51
rect -1 -80 1 -77
rect -1 -91 1 -90
rect -1 -114 1 -111
rect -1 -125 1 -124
<< ndiffusion >>
rect -10 -86 -1 -80
rect -6 -90 -1 -86
rect 1 -84 6 -80
rect 1 -90 10 -84
rect -10 -120 -1 -114
rect -6 -124 -1 -120
rect 1 -118 6 -114
rect 1 -124 10 -118
<< pdiffusion >>
rect -6 26 -1 30
rect -10 6 -1 26
rect 1 6 6 30
rect -6 -31 -1 -27
rect -10 -51 -1 -31
rect 1 -47 10 -27
rect 1 -51 6 -47
<< metal1 >>
rect -21 40 -17 44
rect -13 40 -9 44
rect -5 40 -1 44
rect 3 40 7 44
rect 11 40 15 44
rect -10 30 -6 40
rect -22 1 -3 5
rect 6 -16 10 6
rect -10 -20 10 -16
rect -10 -27 -6 -20
rect -21 -56 -3 -52
rect 6 -68 10 -51
rect 6 -72 28 -68
rect 6 -80 10 -72
rect -10 -103 -6 -90
rect 3 -95 28 -91
rect -10 -107 10 -103
rect 6 -114 10 -107
rect -10 -139 -6 -124
rect 3 -129 15 -125
rect -19 -143 -15 -139
rect -11 -143 -7 -139
rect -3 -143 1 -139
rect 5 -143 9 -139
rect 13 -143 17 -139
<< ntransistor >>
rect -1 -90 1 -80
rect -1 -124 1 -114
<< ptransistor >>
rect -1 6 1 30
rect -1 -51 1 -27
<< polycontact >>
rect -3 1 1 5
rect -3 -56 1 -52
rect -1 -95 3 -91
rect -1 -129 3 -125
<< ndcontact >>
rect -10 -90 -6 -86
rect 6 -84 10 -80
rect -10 -124 -6 -120
rect 6 -118 10 -114
<< pdcontact >>
rect -10 26 -6 30
rect 6 6 10 30
rect -10 -31 -6 -27
rect 6 -51 10 -47
<< psubstratepcontact >>
rect -23 -143 -19 -139
rect -15 -143 -11 -139
rect -7 -143 -3 -139
rect 1 -143 5 -139
rect 9 -143 13 -139
rect 17 -143 21 -139
<< nsubstratencontact >>
rect -25 40 -21 44
rect -17 40 -13 44
rect -9 40 -5 44
rect -1 40 3 44
rect 7 40 11 44
rect 15 40 19 44
<< labels >>
rlabel metal1 -22 1 -22 5 1 vbias1
rlabel metal1 5 42 5 42 1 vdd
rlabel metal1 -21 -56 -21 -52 1 vbias2
rlabel metal1 28 -72 28 -68 7 vout
rlabel metal1 28 -95 28 -91 7 vbias3
rlabel metal1 15 -129 15 -125 1 vin
rlabel metal1 -1 -141 -1 -141 1 gnd
<< end >>
